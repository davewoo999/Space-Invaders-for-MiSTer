//============================================================================
//  Arcade: Space Invaders
//
//  
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//
//  You should have received a copy of the GNU General Public License along
//  with this program; if not, write to the Free Software Foundation, Inc.,
//  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
//============================================================================

// Variuos ports combined -  changes to rom and ram for MiSTer port - Dave Wood (oldgit)
// latest sound module and changes for 2 player added - OSD options to change dip switches

module emu
(
	//Master input clock
	input         CLK_50M,

	//Async reset from top-level module.
	//Can be used as initial reset.
	input         RESET,

	//Must be passed to hps_io module
	inout  [44:0] HPS_BUS,

	//Base video clock. Usually equals to CLK_SYS.
	output        VGA_CLK,

	//Multiple resolutions are supported using different VGA_CE rates.
	//Must be based on CLK_VIDEO
	output        VGA_CE,

	output  [7:0] VGA_R,
	output  [7:0] VGA_G,
	output  [7:0] VGA_B,
	output        VGA_HS,
	output        VGA_VS,
	output        VGA_DE,    // = ~(VBlank | HBlank)

	//Base video clock. Usually equals to CLK_SYS.
	output        HDMI_CLK,

	//Multiple resolutions are supported using different HDMI_CE rates.
	//Must be based on CLK_VIDEO
	output        HDMI_CE,

	output  [7:0] HDMI_R,
	output  [7:0] HDMI_G,
	output  [7:0] HDMI_B,
	output        HDMI_HS,
	output        HDMI_VS,
	output        HDMI_DE,   // = ~(VBlank | HBlank)
	output  [1:0] HDMI_SL,   // scanlines fx

	//Video aspect ratio for HDMI. Most retro systems have ratio 4:3.
	output  [7:0] HDMI_ARX,
	output  [7:0] HDMI_ARY,

	output        LED_USER,  // 1 - ON, 0 - OFF.

	// b[1]: 0 - LED status is system status OR'd with b[0]
	//       1 - LED status is controled solely by b[0]
	// hint: supply 2'b00 to let the system control the LED.
	output  [1:0] LED_POWER,
	output  [1:0] LED_DISK,

	output [15:0] AUDIO_L,
	output [15:0] AUDIO_R,
	output        AUDIO_S    // 1 - signed audio samples, 0 - unsigned
);

assign LED_USER  = ioctl_download;
assign LED_DISK  = 0;
assign LED_POWER = 0;

assign HDMI_ARX = status[1] ? 8'd16 : status[2] ? 8'd4 : 8'd1;
assign HDMI_ARY = status[1] ? 8'd9  : status[2] ? 8'd3 : 8'd1;

`include "build_id.v" 
localparam CONF_STR = {
	"A.invaders;;",
	"-;",
//	"O1,Aspect Ratio,Original,Wide;", --- no effect
//	"O2,Orientation,Vert,Horz;",		 --- cannot get it to work
	"O34,Scanlines(vert),No,25%,50%,75%;",
	"-;",
	"O5,Display Coin Info,ON,OFF;",
//	"O6,Bonus Base,1500pts,1000pts;", This can only be set before game start - changes freezes play and no reset - could add code to reset on change??
	"O78,Bases,3,4,5,6;",
	"-;",
	"-;",
	"T6,Reset;",
	"V,v2.00.",`BUILD_DATE
};

////////////////////   CLOCKS   ///////////////////

wire clk_39p9, clk_9p9, clk_19p9, clk_79p9, clk_4p9;
wire pll_locked;
//wire clk_hdmi;

pll pll
(
	.refclk(CLK_50M),
	.rst(0),
	.outclk_0(clk_79p9),	// 79.870129	x8  79.872
	.outclk_1(clk_39p9),	// 39.935064	x4  39.936
	.outclk_2(clk_19p9),	// 19.967532	x2  19.968
	.outclk_3(clk_9p9),	// 9.983766    should be 9.984 original clk speed
	.outclk_4(clk_4p9),	// 4.991883		/ 2
	.locked(pll_locked)
);


///////////////////////////////////////////////////

wire [31:0] status;
wire  [1:0] buttons;

wire        ioctl_download;
wire        ioctl_wr;
wire [24:0] ioctl_addr;
wire  [7:0] ioctl_dout;

wire [10:0] ps2_key;

wire [15:0] joystick_0, joystick_1;
wire [15:0] joy = joystick_0 | joystick_1;


hps_io #(.STRLEN($size(CONF_STR)>>3)) hps_io
(
	.clk_sys(clk_19p9),
	.HPS_BUS(HPS_BUS),

	.conf_str(CONF_STR),

	.buttons(buttons),
	.status(status),


	.ioctl_download(ioctl_download),
	.ioctl_wr(ioctl_wr),
	.ioctl_addr(ioctl_addr),
	.ioctl_dout(ioctl_dout),

	.joystick_0(joystick_0),
	.joystick_1(joystick_1),
	.ps2_key(ps2_key)
);

wire       pressed = ps2_key[9];
wire [8:0] code    = ps2_key[8:0];
always @(posedge clk_19p9) begin
	reg old_state;
	old_state <= ps2_key[10];
	
	if(old_state != ps2_key[10]) begin
		casex(code)
			'h029: btn_fire         <= pressed; // space
			'h005: btn_one_player   <= pressed; // F1
			'h006: btn_two_players  <= pressed; // F2
			'h01C: btn_left      	<= pressed; // A
			'h023: btn_right      	<= pressed; // D
			'h021: btn_coin  		<= pressed; // C
		endcase
	end
end

reg btn_right = 0;
reg btn_left = 0;
reg btn_one_player = 0;
reg btn_two_players = 0;
reg btn_fire = 0;
reg btn_coin = 0;

wire hblank, vblank;
wire ce_vid = 1; // was clk_9p9
wire hs, vs;
wire rde, rhs, rvs;
wire [2:0] r,g,rr,rg;
wire [2:0] b,rb;

assign VGA_CLK  = clk_19p9; // was clk_19p9
assign VGA_CE   = ce_vid;
//assign VGA_R    = {r,r,r[2:1]};
//assign VGA_G    = {g,g,g[2:1]};
//assign VGA_B    = {b,b,b[2:1]};
//assign VGA_DE   = ~(hblank | vblank);
//assign VGA_HS   = ~hs;
//assign VGA_VS   = ~vs;

assign HDMI_CLK = status[2] ? VGA_CLK: clk_39p9;
assign HDMI_CE  = status[2] ? VGA_CE : 1'b1;
assign HDMI_R   = status[2] ? VGA_R  : {rr,rr,rr[2:1]};
assign HDMI_G   = status[2] ? VGA_G  : {rg,rg,rg[2:1]};
assign HDMI_B   = status[2] ? VGA_B  : {rb,rb,rb[2:1]};
assign HDMI_DE  = status[2] ? VGA_DE : rde;
assign HDMI_HS  = status[2] ? VGA_HS : rhs;
assign HDMI_VS  = status[2] ? VGA_VS : rvs;
assign HDMI_SL  = status[2] ? 2'd0   : status[4:3];

screen_rotate #(318,260,9,2,1,1) screen_rotate
(
	.clk_in(clk_4p9), // with 39.9 hdmi -- 9.9 full height  half width 19.9 double height half width
	.ce_in(ce_vid),
	.video_in({r,g,b}),
	.hblank(hblank),
	.vblank(vblank),

	.clk_out(clk_39p9),
	.video_out({rr,rg,rb}),
	.hsync(rhs),
	.vsync(rvs),
	.de(rde)
);
wire info;
//wire bonus;
wire [1:0] bases;
assign info = status[5];
//assign bonus = status[6];
assign bases = status[8:7];
wire [7:0] audio;
assign AUDIO_L = {audio, audio};
assign AUDIO_R = AUDIO_L;
assign AUDIO_S = 0;

invaders_top invaders_top
(

	.Clk(clk_9p9),
	.Clk_x2(clk_19p9),
	.Clk_x4(clk_39p9),

	.I_RESET(RESET | status[0] | status[6] | buttons[1] | ioctl_download),

	.dn_addr(ioctl_addr[15:0]),
	.dn_data(ioctl_dout),
	.dn_wr(ioctl_wr),

	.video_r(r),
	.video_g(g),
	.video_b(b),
	.video_hblank(hblank),
	.video_vblank(vblank),
	.video_hs(hs),
	.video_vs(vs),
	
	.r(VGA_R),
	.g(VGA_G),
	.b(VGA_B),
	.de(VGA_DE),
	.hs(VGA_HS),
	.vs(VGA_VS),
	
	.audio_out(audio),
	.info(info),
//	.bonus(bonus),
	.bases(bases),
	.btn_coin(btn_coin | joy[8]),
	.btn_one_player(btn_one_player | joy[8]),
	.btn_two_player(btn_two_players),

	.btn_fire(btn_fire | joy[5]),
	.btn_right(btn_right | joy[0]),
	.btn_left(btn_left | joy[1])

);

endmodule
